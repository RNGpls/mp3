library verilog;
use verilog.vl_types.all;
entity zextsh_sv_unit is
end zextsh_sv_unit;
