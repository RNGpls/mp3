library verilog;
use verilog.vl_types.all;
entity byte_extend_sv_unit is
end byte_extend_sv_unit;
